library ieee;
use ieee.std_logic_1164.all;

package components is



end components;